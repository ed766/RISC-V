`include "ALU_TB.sv"
`include "ALU_Control.sv"
`include "CLA_64bit.sv"
`include "Subtractor_64bit.sv"
`include "Array_Multiplier.sv"
`include "abs.sv"