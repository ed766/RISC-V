`include "parameters.sv"
`include "CPU_Core.sv"
`include "ALU.sv"
`include "ALU_Control.sv"
`include "CLA_64bit.sv"
`include "Subtractor_64bit.sv"
`include "Array_Multiplier.sv"
`include "Divider.sv"
`include "register.sv"
